module test();

    if ()
    begin

    end
    else if ()
    begin

    end
        else if ()
        begin

        end
    else
    begin

    end


endmodule
